module main;
initial $runXyceWithDAC;
endmodule

