* Test Netlist
* Simple transient circuit
V1 1 0 SIN(0 1 1)
R1 1 2 50
R2 2 0 100
C1 1 0 1e-6

.TRAN 0 1
.PRINT TRAN V(1) V(2) R1:R TEMP I(V1) I(R1)
.MEASURE TRAN MAXV1 MAX V(1)
.MEASURE TRAN MINV1 MIN V(1)
.MEASURE TRAN MAXV2 MAX V(2)
.MEASURE TRAN MINV2 MIN V(2)


.END

