* a simple high pass filter and low pass filter
*
* high pass cutoff frequency  f = 1/(2 Pi R C)
* R=1000, C=1e-8 f = 16 kHz
* 
* low pass cutoff frequency  f = 1/(2 Pi R C)
* R=1000, C=230e-9 f=690 Hz

* input to filter
ydac dacdriver1 Node1 0 

v1 Node2 0 5.0
v2 Node3 0 -3.0

Ccap Node1 Node2 C=1e-8
Rload Node2 0    R=1000

* output from filter
yadc adchigh Node2 0 simpleADC R=1T
yadc adclow  Node3 0 simpleADC R=1T

* need ref. to ground
rPathToGround1 Node1 0 1e6

rload2 Node1 Node3 R=1000
Clow Node3 0 C=223.0e-9

.model simpleDAC DAC(tr=5e-9 tf=5e-9)
.model simpleADC ADC(settlingtime=5ns uppervoltagelimit=5 lowervoltagelimit=-5)

.print tran V(Node1) v(Node2) v(Node3)
.tran 0 5e-3

.end
