* Test Netlist
* Simple transient circuit
V1 1 0 SIN(0 1 1)
R1 1 0 1
C1 1 0 1e-6

.TRAN 0 1
.PRINT TRAN V(1)
.MEASURE TRAN MAXV1 MAX V(1)
.MEASURE TRAN MINV1 MIN V(1)

.END

