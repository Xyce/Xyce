* Verilog-A vbic_4T_et_cf test circuit
.verilog "vbic_4T_et_cf.vla"

vbe bx 0  0
vcb cx bx 0
vib bx b  0
vic cx c  0
rxth dt 0 1e12
aq1 c  b  0  0 dt vbic
+ RCX=10 RCI=10 RBX=1 RBI=10 RE=1 RBP=10 RS=10
+ IBEN=1.0e-13 RTH=100

.dc vbe 0.5 1.0 0.02
.print dc i(vib) i(vic)
.end
