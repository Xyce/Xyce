module main;
initial $runXyce;
endmodule

