*Sample netlist for BSIM6
*Inverter Transient

*.option abstol=1e-6 reltol=1e-6 post ingold
.options nonlin abstol=1e-6 reltol=1e-6
.options nonlin-tran abstol=1e-6 reltol=1e-6 
.options timeint abstol=1e-6 reltol=1e-6
.options device temp=25

*.hdl "bsim6.va"
.include "modelcard_xyce.nmos"
.include "modelcard_xyce.pmos"

* --- Voltage Sources ---
vdd   supply  0 dc 1.0
vin  vi  0 dc 0.5 sin (0.5 0.5 1MEG)

* --- Inverter Subcircuit ---
.subckt inverter vin vout vdd gnd
Mp1 vout vin vdd gnd pmos W=10u L=10u 
Mn1 vout vin gnd gnd nmos W=10u L=10u 
.ends

* --- Inverter ---
Xinv1  vi 1 supply 0 inverter
Xinv2  1 2 supply 0 inverter
Xinv3  2 3 supply 0 inverter
Xinv4  3 4 supply 0 inverter
Xinv5  4 vo supply 0 inverter

* --- Transient Analysis ---
.tran 10n 5u

.print tran v(vi) v(1) v(2) v(3) v(4) v(vo)

.end
